**Test
.GLOBAL vss! vdd!
.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    HIER_DELIM=0
.options accurate=1 NUMDGT=8 measdgt=5 GMINDC=1e-18 DELMAX=1n method=gear INGOLD=2 POST=1
.INCLUDE "/cae/apps/data/asap7PDK-2022/asap7PDK_r1p7/models/hspice/7nm_TT_160803.pm"
.INCLUDE "MULT2.pex.netlist"

**Set up power rails
v1 vdd! 0 0.9v
v2 vss! 0 0v

**Stimulus
v3 A 0 pwl 	0ns 0.9v  2ns 0.9v  2.025ns 0v  9ns 0v 
v4 B 0 pwl 	0ns 0.9v  3ns 0.9v  3.025ns 0v  6ns 0v  6.025ns 0.9v  9ns 0.9v 
v5 Cin 0 pwl 	0ns 0.9v 

X_DUT vss! vdd! B<1> A<1> B<0> A<0> out_Y<0> out_Y<1> CONVFA

.OP
.TRAN STEP=10p STOP=9n
.end
