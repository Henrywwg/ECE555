* SPICE NETLIST
***************************************

.SUBCKT neuron vss vdd w0<1> x0<1> w0<0> x0<0> w1<0> x1<0> w1<1> x1<1> w2<0> w2<1> w2<2> Z<2> Z<0> Z<1>
** N=538 EP=16 IP=0 FDC=326
M0 5 w0<1> vss vss nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-8572 $Y=4428 $D=1
M1 6 x0<1> vss vss nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-8572 $Y=6048 $D=1
M2 80 5 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-7924 $Y=4428 $D=1
M3 81 6 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-7924 $Y=6156 $D=1
M4 12 x0<1> 80 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-7708 $Y=4428 $D=1
M5 14 w0<1> 81 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-7708 $Y=6156 $D=1
M6 82 5 12 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-7492 $Y=4428 $D=1
M7 83 6 14 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-7492 $Y=6156 $D=1
M8 vss x0<1> 82 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-7276 $Y=4428 $D=1
M9 vss w0<1> 83 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-7276 $Y=6156 $D=1
M10 84 7 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6628 $Y=108 $D=1
M11 29 9 72 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6628 $Y=1836 $D=1
M12 85 8 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6628 $Y=2268 $D=1
M13 18 10 84 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6412 $Y=108 $D=1
M14 72 9 29 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6412 $Y=1836 $D=1
M15 15 11 85 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6412 $Y=2268 $D=1
M16 86 8 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6412 $Y=3996 $D=1
M17 87 12 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6412 $Y=4428 $D=1
M18 88 w0<0> vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6412 $Y=6048 $D=1
M19 89 7 18 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6196 $Y=108 $D=1
M20 90 8 15 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6196 $Y=2268 $D=1
M21 21 15 86 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6196 $Y=3996 $D=1
M22 22 14 87 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6196 $Y=4428 $D=1
M23 17 x0<0> 88 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-6196 $Y=6048 $D=1
M24 vss 10 89 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5980 $Y=108 $D=1
M25 vss 11 90 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5980 $Y=2268 $D=1
M26 91 8 21 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5980 $Y=3996 $D=1
M27 92 12 22 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5980 $Y=4428 $D=1
M28 93 x0<0> 17 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5980 $Y=6048 $D=1
M29 72 8 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5764 $Y=1836 $D=1
M30 vss 15 91 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5764 $Y=3996 $D=1
M31 vss 14 92 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5764 $Y=4428 $D=1
M32 vss w0<0> 93 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5764 $Y=6048 $D=1
M33 vss 11 72 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5548 $Y=1836 $D=1
M34 10 17 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5548 $Y=6048 $D=1
M35 33 18 73 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5332 $Y=108 $D=1
M36 72 11 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5332 $Y=1836 $D=1
M37 73 18 33 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5116 $Y=108 $D=1
M38 vss 8 72 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5116 $Y=1836 $D=1
M39 94 15 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-5116 $Y=2268 $D=1
M40 19 11 94 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4900 $Y=2268 $D=1
M41 95 19 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4900 $Y=3996 $D=1
M42 96 10 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4900 $Y=4536 $D=1
M43 vss 20 8 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4900 $Y=6048 $D=1
M44 97 15 19 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4684 $Y=2268 $D=1
M45 25 21 95 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4684 $Y=3996 $D=1
M46 24 22 96 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4684 $Y=4536 $D=1
M47 98 7 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4684 $Y=6048 $D=1
M48 73 7 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4468 $Y=108 $D=1
M49 99 8 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4468 $Y=1836 $D=1
M50 vss 11 97 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4468 $Y=2268 $D=1
M51 100 19 25 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4468 $Y=3996 $D=1
M52 101 22 24 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4468 $Y=4536 $D=1
M53 20 23 98 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4468 $Y=6048 $D=1
M54 vss 10 73 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4252 $Y=108 $D=1
M55 29 11 99 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4252 $Y=1836 $D=1
M56 vss 21 100 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4252 $Y=3996 $D=1
M57 vss 10 101 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4252 $Y=4536 $D=1
M58 102 23 20 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4252 $Y=6048 $D=1
M59 73 10 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4036 $Y=108 $D=1
M60 103 11 29 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4036 $Y=1836 $D=1
M61 11 24 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4036 $Y=4536 $D=1
M62 vss 7 102 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-4036 $Y=6048 $D=1
M63 vss 7 73 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-3820 $Y=108 $D=1
M64 vss 8 103 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-3820 $Y=1836 $D=1
M65 104 9 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-3604 $Y=2268 $D=1
M66 27 25 104 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-3388 $Y=2268 $D=1
M67 105 9 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-3388 $Y=3996 $D=1
M68 vss 26 7 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-3388 $Y=4536 $D=1
M69 9 18 vss vss nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-3172 $Y=108 $D=1
M70 46 29 vss vss nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-3172 $Y=1728 $D=1
M71 106 9 27 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-3172 $Y=2268 $D=1
M72 35 27 105 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-3172 $Y=3996 $D=1
M73 107 w1<0> vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-3172 $Y=4536 $D=1
M74 108 28 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-3172 $Y=6156 $D=1
M75 vss 25 106 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-2956 $Y=2268 $D=1
M76 109 9 35 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-2956 $Y=3996 $D=1
M77 26 x1<0> 107 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-2956 $Y=4536 $D=1
M78 23 31 108 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-2956 $Y=6156 $D=1
M79 vss 27 109 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-2740 $Y=3996 $D=1
M80 110 x1<0> 26 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-2740 $Y=4536 $D=1
M81 111 28 23 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-2740 $Y=6156 $D=1
M82 44 33 vss vss nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-2524 $Y=108 $D=1
M83 vss w1<0> 110 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-2524 $Y=4536 $D=1
M84 vss 31 111 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-2524 $Y=6156 $D=1
M85 112 27 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-2092 $Y=2268 $D=1
M86 34 25 112 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1876 $Y=2268 $D=1
M87 113 34 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1876 $Y=3996 $D=1
M88 114 27 34 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1660 $Y=2268 $D=1
M89 45 35 113 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1660 $Y=3996 $D=1
M90 115 w1<1> vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1660 $Y=4428 $D=1
M91 116 x1<1> vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1660 $Y=6156 $D=1
M92 vss 25 114 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1444 $Y=2268 $D=1
M93 117 34 45 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1444 $Y=3996 $D=1
M94 28 38 115 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1444 $Y=4428 $D=1
M95 31 39 116 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1444 $Y=6156 $D=1
M96 vss 35 117 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1228 $Y=3996 $D=1
M97 118 w1<1> 28 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1228 $Y=4428 $D=1
M98 119 x1<1> 31 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1228 $Y=6156 $D=1
M99 vss 38 118 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1012 $Y=4428 $D=1
M100 vss 39 119 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=-1012 $Y=6156 $D=1
M101 vss x1<1> 38 vss nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-364 $Y=4428 $D=1
M102 vss w1<1> 39 vss nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-364 $Y=6048 $D=1
M103 120 w2<0> vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=284 $Y=108 $D=1
M104 59 43 75 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=284 $Y=1836 $D=1
M105 121 w2<1> vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=284 $Y=2268 $D=1
M106 122 w2<2> vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=284 $Y=4428 $D=1
M107 49 44 120 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=500 $Y=108 $D=1
M108 75 43 59 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=500 $Y=1836 $D=1
M109 47 45 121 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=500 $Y=2268 $D=1
M110 123 w2<1> vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=500 $Y=3996 $D=1
M111 48 46 122 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=500 $Y=4428 $D=1
M112 124 w2<2> vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=500 $Y=6156 $D=1
M113 125 w2<0> 49 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=716 $Y=108 $D=1
M114 126 w2<1> 47 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=716 $Y=2268 $D=1
M115 52 47 123 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=716 $Y=3996 $D=1
M116 127 w2<2> 48 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=716 $Y=4428 $D=1
M117 53 48 124 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=716 $Y=6156 $D=1
M118 vss 44 125 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=932 $Y=108 $D=1
M119 vss 45 126 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=932 $Y=2268 $D=1
M120 128 w2<1> 52 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=932 $Y=3996 $D=1
M121 vss 46 127 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=932 $Y=4428 $D=1
M122 129 w2<2> 53 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=932 $Y=6156 $D=1
M123 75 w2<1> vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1148 $Y=1836 $D=1
M124 vss 47 128 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1148 $Y=3996 $D=1
M125 vss 48 129 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1148 $Y=6156 $D=1
M126 vss 45 75 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1364 $Y=1836 $D=1
M127 60 49 76 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1580 $Y=108 $D=1
M128 75 45 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1580 $Y=1836 $D=1
M129 76 49 60 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1796 $Y=108 $D=1
M130 vss w2<1> 75 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1796 $Y=1836 $D=1
M131 130 47 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1796 $Y=2268 $D=1
M132 131 48 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=1796 $Y=4428 $D=1
M133 50 45 130 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2012 $Y=2268 $D=1
M134 132 50 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2012 $Y=3996 $D=1
M135 51 46 131 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2012 $Y=4428 $D=1
M136 133 51 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2012 $Y=6156 $D=1
M137 134 47 50 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2228 $Y=2268 $D=1
M138 55 52 132 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2228 $Y=3996 $D=1
M139 135 48 51 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2228 $Y=4428 $D=1
M140 56 53 133 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2228 $Y=6156 $D=1
M141 76 w2<0> vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2444 $Y=108 $D=1
M142 136 w2<1> vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2444 $Y=1836 $D=1
M143 vss 45 134 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2444 $Y=2268 $D=1
M144 137 50 55 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2444 $Y=3996 $D=1
M145 vss 46 135 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2444 $Y=4428 $D=1
M146 138 51 56 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2444 $Y=6156 $D=1
M147 vss 44 76 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2660 $Y=108 $D=1
M148 59 45 136 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2660 $Y=1836 $D=1
M149 vss 52 137 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2660 $Y=3996 $D=1
M150 vss 53 138 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2660 $Y=6156 $D=1
M151 76 44 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2876 $Y=108 $D=1
M152 139 45 59 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=2876 $Y=1836 $D=1
M153 vss w2<0> 76 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3092 $Y=108 $D=1
M154 vss w2<1> 139 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3092 $Y=1836 $D=1
M155 140 43 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3308 $Y=2268 $D=1
M156 141 54 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3308 $Y=4428 $D=1
M157 57 55 140 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3524 $Y=2268 $D=1
M158 142 43 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3524 $Y=3996 $D=1
M159 58 56 141 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3524 $Y=4428 $D=1
M160 143 54 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3524 $Y=6156 $D=1
M161 43 49 vss vss nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3740 $Y=108 $D=1
M162 54 59 vss vss nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3740 $Y=1728 $D=1
M163 144 43 57 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3740 $Y=2268 $D=1
M164 63 57 142 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3740 $Y=3996 $D=1
M165 145 54 58 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3740 $Y=4428 $D=1
M166 64 58 143 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3740 $Y=6156 $D=1
M167 vss 55 144 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3956 $Y=2268 $D=1
M168 146 43 63 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3956 $Y=3996 $D=1
M169 vss 56 145 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3956 $Y=4428 $D=1
M170 147 54 64 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=3956 $Y=6156 $D=1
M171 vss 57 146 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4172 $Y=3996 $D=1
M172 vss 58 147 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4172 $Y=6156 $D=1
M173 65 60 vss vss nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4388 $Y=108 $D=1
M174 148 57 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4820 $Y=2268 $D=1
M175 149 58 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=4820 $Y=4428 $D=1
M176 61 55 148 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5036 $Y=2268 $D=1
M177 150 61 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5036 $Y=3996 $D=1
M178 62 56 149 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5036 $Y=4428 $D=1
M179 151 62 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5036 $Y=6156 $D=1
M180 152 57 61 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5252 $Y=2268 $D=1
M181 66 63 150 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5252 $Y=3996 $D=1
M182 153 58 62 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5252 $Y=4428 $D=1
M183 67 64 151 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5252 $Y=6156 $D=1
M184 vss 55 152 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5468 $Y=2268 $D=1
M185 154 61 66 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5468 $Y=3996 $D=1
M186 vss 56 153 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5468 $Y=4428 $D=1
M187 155 62 67 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5468 $Y=6156 $D=1
M188 vss 63 154 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5684 $Y=3996 $D=1
M189 vss 64 155 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=5684 $Y=6156 $D=1
M190 156 65 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=6332 $Y=2376 $D=1
M191 157 66 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=6332 $Y=3888 $D=1
M192 68 67 vss vss nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6332 $Y=4428 $D=1
M193 69 68 156 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=6548 $Y=2376 $D=1
M194 70 68 157 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=6548 $Y=3888 $D=1
M195 158 68 69 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=6764 $Y=2376 $D=1
M196 159 68 70 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=6764 $Y=3888 $D=1
M197 vss 65 158 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=6980 $Y=2376 $D=1
M198 vss 66 159 vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=6980 $Y=3888 $D=1
M199 Z<0> 69 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7196 $Y=2376 $D=1
M200 Z<1> 70 vss vss nmos_rvt L=2e-08 W=5.4e-08 nfin=2 $X=7196 $Y=3888 $D=1
M201 Z<2> vdd vss vss nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7196 $Y=4428 $D=1
M202 5 w0<1> vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-8572 $Y=4968 $D=0
M203 6 x0<1> vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-8572 $Y=5508 $D=0
M204 12 x0<1> vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-7708 $Y=4968 $D=0
M205 14 w0<1> vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-7708 $Y=5508 $D=0
M206 vdd 5 12 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-7492 $Y=4968 $D=0
M207 vdd 6 14 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-7492 $Y=5508 $D=0
M208 29 9 71 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-6628 $Y=1188 $D=0
M209 18 10 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-6412 $Y=648 $D=0
M210 71 9 29 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-6412 $Y=1188 $D=0
M211 15 11 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-6412 $Y=2808 $D=0
M212 17 w0<0> vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-6412 $Y=5508 $D=0
M213 vdd 7 18 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-6196 $Y=648 $D=0
M214 vdd 8 15 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-6196 $Y=2808 $D=0
M215 21 15 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-6196 $Y=3348 $D=0
M216 22 14 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-6196 $Y=4968 $D=0
M217 vdd x0<0> 17 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-6196 $Y=5508 $D=0
M218 vdd 8 21 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-5980 $Y=3348 $D=0
M219 vdd 12 22 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-5980 $Y=4968 $D=0
M220 71 8 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-5764 $Y=1188 $D=0
M221 vdd 11 71 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-5548 $Y=1188 $D=0
M222 10 17 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-5548 $Y=5508 $D=0
M223 33 18 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-5332 $Y=648 $D=0
M224 71 11 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-5332 $Y=1188 $D=0
M225 vdd 8 71 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-5116 $Y=1188 $D=0
M226 19 11 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4900 $Y=2808 $D=0
M227 24 10 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4900 $Y=4968 $D=0
M228 vdd 20 8 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4900 $Y=5508 $D=0
M229 vdd 15 19 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4684 $Y=2808 $D=0
M230 25 21 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4684 $Y=3348 $D=0
M231 vdd 22 24 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4684 $Y=4968 $D=0
M232 160 7 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4468 $Y=648 $D=0
M233 161 8 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4468 $Y=1188 $D=0
M234 vdd 19 25 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4468 $Y=3348 $D=0
M235 33 10 160 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4252 $Y=648 $D=0
M236 29 11 161 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4252 $Y=1188 $D=0
M237 20 23 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4252 $Y=5508 $D=0
M238 162 10 33 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4036 $Y=648 $D=0
M239 163 11 29 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4036 $Y=1188 $D=0
M240 11 24 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4036 $Y=4968 $D=0
M241 vdd 7 20 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-4036 $Y=5508 $D=0
M242 vdd 7 162 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-3820 $Y=648 $D=0
M243 vdd 8 163 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-3820 $Y=1188 $D=0
M244 27 25 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-3388 $Y=2808 $D=0
M245 vdd 26 7 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-3388 $Y=4968 $D=0
M246 9 18 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-3172 $Y=648 $D=0
M247 46 29 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-3172 $Y=1188 $D=0
M248 vdd 9 27 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-3172 $Y=2808 $D=0
M249 35 27 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-3172 $Y=3348 $D=0
M250 vdd 9 35 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-2956 $Y=3348 $D=0
M251 23 31 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-2956 $Y=5508 $D=0
M252 26 x1<0> vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-2740 $Y=4968 $D=0
M253 vdd 28 23 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-2740 $Y=5508 $D=0
M254 44 33 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-2524 $Y=648 $D=0
M255 vdd w1<0> 26 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-2524 $Y=4968 $D=0
M256 34 25 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-1876 $Y=2808 $D=0
M257 vdd 27 34 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-1660 $Y=2808 $D=0
M258 45 35 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-1660 $Y=3348 $D=0
M259 vdd 34 45 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-1444 $Y=3348 $D=0
M260 28 38 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-1444 $Y=4968 $D=0
M261 31 39 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-1444 $Y=5508 $D=0
M262 vdd w1<1> 28 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-1228 $Y=4968 $D=0
M263 vdd x1<1> 31 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-1228 $Y=5508 $D=0
M264 vdd x1<1> 38 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-364 $Y=4968 $D=0
M265 vdd w1<1> 39 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=-364 $Y=5508 $D=0
M266 59 43 74 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=284 $Y=1188 $D=0
M267 49 44 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=500 $Y=648 $D=0
M268 74 43 59 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=500 $Y=1188 $D=0
M269 47 45 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=500 $Y=2808 $D=0
M270 48 46 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=500 $Y=4968 $D=0
M271 vdd w2<0> 49 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=716 $Y=648 $D=0
M272 vdd w2<1> 47 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=716 $Y=2808 $D=0
M273 52 47 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=716 $Y=3348 $D=0
M274 vdd w2<2> 48 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=716 $Y=4968 $D=0
M275 53 48 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=716 $Y=5508 $D=0
M276 vdd w2<1> 52 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=932 $Y=3348 $D=0
M277 vdd w2<2> 53 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=932 $Y=5508 $D=0
M278 74 w2<1> vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1148 $Y=1188 $D=0
M279 vdd 45 74 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1364 $Y=1188 $D=0
M280 60 49 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1580 $Y=648 $D=0
M281 74 45 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1580 $Y=1188 $D=0
M282 vdd w2<1> 74 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=1796 $Y=1188 $D=0
M283 50 45 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2012 $Y=2808 $D=0
M284 51 46 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2012 $Y=4968 $D=0
M285 vdd 47 50 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2228 $Y=2808 $D=0
M286 55 52 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2228 $Y=3348 $D=0
M287 vdd 48 51 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2228 $Y=4968 $D=0
M288 56 53 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2228 $Y=5508 $D=0
M289 164 w2<0> vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2444 $Y=648 $D=0
M290 165 w2<1> vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2444 $Y=1188 $D=0
M291 vdd 50 55 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2444 $Y=3348 $D=0
M292 vdd 51 56 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2444 $Y=5508 $D=0
M293 60 44 164 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2660 $Y=648 $D=0
M294 59 45 165 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2660 $Y=1188 $D=0
M295 166 44 60 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2876 $Y=648 $D=0
M296 167 45 59 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=2876 $Y=1188 $D=0
M297 vdd w2<0> 166 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3092 $Y=648 $D=0
M298 vdd w2<1> 167 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3092 $Y=1188 $D=0
M299 57 55 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3524 $Y=2808 $D=0
M300 58 56 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3524 $Y=4968 $D=0
M301 43 49 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3740 $Y=648 $D=0
M302 54 59 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3740 $Y=1188 $D=0
M303 vdd 43 57 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3740 $Y=2808 $D=0
M304 63 57 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3740 $Y=3348 $D=0
M305 vdd 54 58 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3740 $Y=4968 $D=0
M306 64 58 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3740 $Y=5508 $D=0
M307 vdd 43 63 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3956 $Y=3348 $D=0
M308 vdd 54 64 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=3956 $Y=5508 $D=0
M309 65 60 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=4388 $Y=648 $D=0
M310 61 55 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5036 $Y=2808 $D=0
M311 62 56 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5036 $Y=4968 $D=0
M312 vdd 57 61 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5252 $Y=2808 $D=0
M313 66 63 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5252 $Y=3348 $D=0
M314 vdd 58 62 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5252 $Y=4968 $D=0
M315 67 64 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5252 $Y=5508 $D=0
M316 vdd 61 66 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5468 $Y=3348 $D=0
M317 vdd 62 67 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=5468 $Y=5508 $D=0
M318 69 65 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6332 $Y=2808 $D=0
M319 70 66 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6332 $Y=3348 $D=0
M320 68 67 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6332 $Y=4968 $D=0
M321 vdd 68 69 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6548 $Y=2808 $D=0
M322 vdd 68 70 vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=6548 $Y=3348 $D=0
M323 Z<0> 69 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7196 $Y=2808 $D=0
M324 Z<1> 70 vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7196 $Y=3348 $D=0
M325 Z<2> vdd vdd vdd pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=7196 $Y=4968 $D=0
.ENDS
***************************************
